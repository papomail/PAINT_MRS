�� z  �   �zHa=1���y�a=1�� gamma 1�{K)���z�)�� gamma 2��4�̣���̣ alpha 1��u��v���C��v� alpha 2���!(�;����!(�;� beta 1��kn�O����Rn�O�� beta 2����S.{>����S.{> beta 3��d���vB��2���vB NAD        @)       PCr@}P�:h��@~�:h�� GPC@���+�D@��+�D GPE@�!�����@������� Pi@��Cϳ1@�Cϳ1 Pi_2@��0U2a@�@�0U2a PME@�Fky��@�xky�� PCh��O�X������X��� UDP@�@?���@��?��� Pi_3@�S��%��@����%�� PME2@���A_E�@��A_E� Pi4