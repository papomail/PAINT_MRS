�� z     @���c�A @�H�c�A  Naa_2CH3@��=� �@�"=� � Cho@�
8���@�28��� GPC@���J���@��J��� 	Cr_N(CH3)@�X�{9@���{9 Cr_2CH2@�X���c@�����c NaaG@�;Q�\л@��Q�\л Lac1@�[Ho��V@��Ho��V Lac2@�ٲ�s�@���s� Glycine@��Ğ�z@�@Ğ�z Al1@�6�����@������� Al2