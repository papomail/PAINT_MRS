�� w�   ����d���#��r�8� w1@,��P��S@E�=<b�_ w2�,��P���@���5 w3�{�m�n��|�DR�&� F1�}�4)�:�����r� F2�v�]�	�tkb��{ F3