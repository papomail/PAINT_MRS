�� z  �   �`ͣ�,�#�^{G�Y�F gamma 1�asc�_�_�,�",� gamma 2�x��(��w��(� alpha 1�x�^�A�x�^�A alpha 2��n�mNs��
�mNs beta 1��i6V���i6V beta 2������f���]���f� beta 3�z�dq ��yK�dq � NAD        @)       PCr@b���Yv�@dM��Yv� GPC@f���-
@h��-
 GPE@p�җDEM@q|җDEM Pi@o�dH<�W@p�2$h, Pi_2@u���u[�@v���u[� PME@t�jXf�@u�jXf� PCh���v��~N��v� UDP@m��� ��@oJ�� �� Pi_3@scn5��@t+n5�� PME2@k�@�&@mZ@�& Pi4